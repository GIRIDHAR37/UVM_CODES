typedef uvm_sequencer#(fifo_wtx) fifo_wsqr;

/*class fifo_wsqr extends uvm_sequencer#(fifo_wtx);
	
	`uvm_component_utils(fifo_wsqr)

	function new(string name="",uvm_component parent);
		super.new(name,parent);
	endfunction

	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
	endfunction

endclass*/
