interface lg_if();
	logic [3:0]a;
	logic [3:0]b;
	logic [2:0]mode;
	logic [3:0]y;
endinterface

