interface pd_if(input bit clk,rst);
	logic data;
	logic valid;
	logic pd_o;
endinterface
