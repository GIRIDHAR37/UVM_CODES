typedef uvm_sequencer#(fifo_tx) fifo_sqr;

/*class fifo_sqr extends uvm_sequencer#(fifo_tx);
	
	`uvm_component_utils(fifo_sqr)

	function new(string name="",uvm_component parent);
		super.new(name,parent);
	endfunction

	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
	endfunction

endclass*/
