typedef uvm_sequencer#(fifo_rtx) fifo_rsqr;

/*class fifo_rsqr extends uvm_sequencer#(fifo_rtx);
	
	`uvm_component_utils(fifo_rsqr)

	function new(string name="",uvm_component parent);
		super.new(name,parent);
	endfunction

	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
	endfunction

endclass*/

